`timescale 1ns / 1ps
`default_nettype none
/***********************************************************************************************************************
*                                                                                                                      *
* ANTIKERNEL                                                                                                           *
*                                                                                                                      *
* Copyright (c) 2012-2024 Andrew D. Zonenberg                                                                          *
* All rights reserved.                                                                                                 *
*                                                                                                                      *
* Redistribution and use in source and binary forms, with or without modification, are permitted provided that the     *
* following conditions are met:                                                                                        *
*                                                                                                                      *
*    * Redistributions of source code must retain the above copyright notice, this list of conditions, and the         *
*      following disclaimer.                                                                                           *
*                                                                                                                      *
*    * Redistributions in binary form must reproduce the above copyright notice, this list of conditions and the       *
*      following disclaimer in the documentation and/or other materials provided with the distribution.                *
*                                                                                                                      *
*    * Neither the name of the author nor the names of any contributors may be used to endorse or promote products     *
*      derived from this software without specific prior written permission.                                           *
*                                                                                                                      *
* THIS SOFTWARE IS PROVIDED BY THE AUTHORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED   *
* TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL *
* THE AUTHORS BE HELD LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES        *
* (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR       *
* BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT *
* (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE       *
* POSSIBILITY OF SUCH DAMAGE.                                                                                          *
*                                                                                                                      *
***********************************************************************************************************************/

`include "GmiiBus.svh"
`include "EthernetBus.svh"

/**
	@file
	@author Andrew D. Zonenberg
	@brief Convenience wrapper around XGEthernetMAC and XGEthernetPCS
 */
module XGMACWrapper(
	//Clocks for transmit/receive domains, generated by the transceiver
	//Both are nominally 312.5 MHz, but may have a slight phase difference
	input wire								rx_clk,
	input wire								tx_clk,

	//Incoming data from the GT's 64/66b gearbox
	input wire								rx_data_valid,
	input wire								rx_header_valid,
	input wire[1:0]							rx_header,
	input wire[31:0]						rx_data,
	output wire								rx_bitslip,

	//Outbound data to the GT's 64/66b gearbox
	output wire[5:0]						tx_sequence,
	output wire[1:0]						tx_header,
	output wire[31:0]						tx_data,

	//Link state etc signals
	input wire								sfp_los,

	//MAC signals to TCP/IP stack
	output wire								mac_rx_clk,
	output EthernetRxBus					mac_rx_bus,

	//note that unlike most 1G variants, TX clock is different from RX
	output wire								mac_tx_clk,
	input wire EthernetTxBus				mac_tx_bus,

	//mac_rx_clk domain
	output wire								link_up,
	//no link speed since we're not dynamic 1G/10G, we only support 10G

	//TODO: performance counters
	output wire								remote_fault
	);

	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// PCS

	assign mac_rx_clk = rx_clk;
	assign mac_tx_clk = tx_clk;

	XgmiiBus xgmii_rx_bus;
	XgmiiBus xgmii_tx_bus;

	XGEthernetPCS pcs(
		.rx_clk(rx_clk),
		.tx_clk(tx_clk),

		.rx_data_valid(rx_data_valid),
		.rx_header_valid(rx_header_valid),
		.rx_header(rx_header),
		.rx_data(rx_data),
		.rx_bitslip(rx_bitslip),

		.tx_sequence(tx_sequence),
		.tx_header(tx_header),
		.tx_data(tx_data),

		.xgmii_rx_clk(),
		.xgmii_rx_bus(xgmii_rx_bus),

		.xgmii_tx_clk(),
		.xgmii_tx_bus(xgmii_tx_bus),

		.sfp_los(sfp_los),
		.block_sync_good(),
		.link_up(link_up),
		.remote_fault(remote_fault)
	);

	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Pipeline register on the XGMII RX bus to improve timing
	// (tight on Kintex7 -2, might be able to remove on ultrascale?)

	XgmiiBus	xgmii_rx_bus_ff;
	always_ff @(posedge mac_rx_clk) begin
		xgmii_rx_bus_ff	<= xgmii_rx_bus;
	end

	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// The actual MAC

	XGEthernetMAC mac(
		.xgmii_rx_clk(mac_rx_clk),
		.xgmii_rx_bus(xgmii_rx_bus_ff),

		.xgmii_tx_clk(mac_tx_clk),
		.xgmii_tx_bus(xgmii_tx_bus),

		.link_up(link_up),

		.rx_bus(mac_rx_bus),
		.tx_bus(mac_tx_bus)

		//TODO: performance counters
	);

endmodule
