`timescale 1ns / 1ps
`default_nettype none
/***********************************************************************************************************************
*                                                                                                                      *
* ANTIKERNEL                                                                                                           *
*                                                                                                                      *
* Copyright (c) 2012-2025 Andrew D. Zonenberg                                                                          *
* All rights reserved.                                                                                                 *
*                                                                                                                      *
* Redistribution and use in source and binary forms, with or without modification, are permitted provided that the     *
* following conditions are met:                                                                                        *
*                                                                                                                      *
*    * Redistributions of source code must retain the above copyright notice, this list of conditions, and the         *
*      following disclaimer.                                                                                           *
*                                                                                                                      *
*    * Redistributions in binary form must reproduce the above copyright notice, this list of conditions and the       *
*      following disclaimer in the documentation and/or other materials provided with the distribution.                *
*                                                                                                                      *
*    * Neither the name of the author nor the names of any contributors may be used to endorse or promote products     *
*      derived from this software without specific prior written permission.                                           *
*                                                                                                                      *
* THIS SOFTWARE IS PROVIDED BY THE AUTHORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED   *
* TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL *
* THE AUTHORS BE HELD LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES        *
* (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR       *
* BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT *
* (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE       *
* POSSIBILITY OF SUCH DAMAGE.                                                                                          *
*                                                                                                                      *
***********************************************************************************************************************/

module GTYLane_UltraScale #(
	parameter FOO = "BAR"
) (

	//APB to DRP
	//DRP space is mapped as 32-bit words with the high 16 bits write-ignored / RAZ
	//Accesses must be aligned
	APB.completer 		apb
);

	GTYE4_CHANNEL #(
		.ACJTAG_DEBUG_MODE(),
		.ACJTAG_MODE(),
		.ACJTAG_RESET(),
		.ADAPT_CFG0(),
		.ADAPT_CFG1(),
		.ADAPT_CFG2(),
		.ALIGN_COMMA_DOUBLE(),
		.ALIGN_COMMA_ENABLE(),
		.ALIGN_COMMA_WORD(),
		.ALIGN_MCOMMA_DET(),
		.ALIGN_MCOMMA_VALUE(),
		.ALIGN_PCOMMA_DET(),
		.ALIGN_PCOMMA_VALUE(),
		.A_RXOSCALRESET(),
		.A_RXPROGDIVRESET(),
		.A_RXTERMINATION(),
		.A_TXDIFFCTRL(),
		.A_TXPROGDIVRESET(),
		.CBCC_DATA_SOURCE_SEL(),
		.CDR_SWAP_MODE_EN(),
		.CFOK_PWRSVE_EN(),
		.CHAN_BOND_KEEP_ALIGN(),
		.CHAN_BOND_MAX_SKEW(),
		.CHAN_BOND_SEQ_1_1(),
		.CHAN_BOND_SEQ_1_2(),
		.CHAN_BOND_SEQ_1_3(),
		.CHAN_BOND_SEQ_1_4(),
		.CHAN_BOND_SEQ_1_ENABLE(),
		.CHAN_BOND_SEQ_2_1(),
		.CHAN_BOND_SEQ_2_2(),
		.CHAN_BOND_SEQ_2_3(),
		.CHAN_BOND_SEQ_2_4(),
		.CHAN_BOND_SEQ_2_ENABLE(),
		.CHAN_BOND_SEQ_2_USE(),
		.CHAN_BOND_SEQ_LEN(),
		.CH_HSPMUX(),
		.CKCAL1_CFG_0(),
		.CKCAL1_CFG_1(),
		.CKCAL1_CFG_2(),
		.CKCAL1_CFG_3(),
		.CKCAL2_CFG_0(),
		.CKCAL2_CFG_1(),
		.CKCAL2_CFG_2(),
		.CKCAL2_CFG_3(),
		.CKCAL2_CFG_4(),
		.CLK_CORRECT_USE(),
		.CLK_COR_KEEP_IDLE(),
		.CLK_COR_MAX_LAT(),
		.CLK_COR_MIN_LAT(),
		.CLK_COR_PRECEDENCE(),
		.CLK_COR_REPEAT_WAIT(),
		.CLK_COR_SEQ_1_1(),
		.CLK_COR_SEQ_1_2(),
		.CLK_COR_SEQ_1_3(),
		.CLK_COR_SEQ_1_4(),
		.CLK_COR_SEQ_1_ENABLE(),
		.CLK_COR_SEQ_2_1(),
		.CLK_COR_SEQ_2_2(),
		.CLK_COR_SEQ_2_3(),
		.CLK_COR_SEQ_2_4(),
		.CLK_COR_SEQ_2_ENABLE(),
		.CLK_COR_SEQ_2_USE(),
		.CLK_COR_SEQ_LEN(),
		.CPLL_CFG0(),
		.CPLL_CFG1(),
		.CPLL_CFG2(),
		.CPLL_CFG3(),
		.CPLL_FBDIV(),
		.CPLL_FBDIV_45(),
		.CPLL_INIT_CFG0(),
		.CPLL_LOCK_CFG(),
		.CPLL_REFCLK_DIV(),
		.CTLE3_OCAP_EXT_CTRL(),
		.CTLE3_OCAP_EXT_EN(),
		.DDI_CTRL(),
		.DDI_REALIGN_WAIT(),
		.DEC_MCOMMA_DETECT(),
		.DEC_PCOMMA_DETECT(),
		.DEC_VALID_COMMA_ONLY(),
		.DELAY_ELEC(),
		.DMONITOR_CFG0(),
		.DMONITOR_CFG1(),
		.ES_CLK_PHASE_SEL(),
		.ES_CONTROL(),
		.ES_ERRDET_EN(),
		.ES_EYE_SCAN_EN(),
		.ES_HORZ_OFFSET(),
		.ES_PRESCALE(),
		.ES_QUALIFIER0(),
		.ES_QUALIFIER1(),
		.ES_QUALIFIER2(),
		.ES_QUALIFIER3(),
		.ES_QUALIFIER4(),
		.ES_QUALIFIER5(),
		.ES_QUALIFIER6(),
		.ES_QUALIFIER7(),
		.ES_QUALIFIER8(),
		.ES_QUALIFIER9(),
		.ES_QUAL_MASK0(),
		.ES_QUAL_MASK1(),
		.ES_QUAL_MASK2(),
		.ES_QUAL_MASK3(),
		.ES_QUAL_MASK4(),
		.ES_QUAL_MASK5(),
		.ES_QUAL_MASK6(),
		.ES_QUAL_MASK7(),
		.ES_QUAL_MASK8(),
		.ES_QUAL_MASK9(),
		.ES_SDATA_MASK0(),
		.ES_SDATA_MASK1(),
		.ES_SDATA_MASK2(),
		.ES_SDATA_MASK3(),
		.ES_SDATA_MASK4(),
		.ES_SDATA_MASK5(),
		.ES_SDATA_MASK6(),
		.ES_SDATA_MASK7(),
		.ES_SDATA_MASK8(),
		.ES_SDATA_MASK9(),
		.EYESCAN_VP_RANGE(),
		.EYE_SCAN_SWAP_EN(),
		.FTS_DESKEW_SEQ_ENABLE(),
		.FTS_LANE_DESKEW_CFG(),
		.FTS_LANE_DESKEW_EN(),
		.GEARBOX_MODE(),
		.ISCAN_CK_PH_SEL2(),
		.LOCAL_MASTER(),
		.LPBK_BIAS_CTRL(),
		.LPBK_EN_RCAL_B(),
		.LPBK_EXT_RCAL(),
		.LPBK_IND_CTRL0(),
		.LPBK_IND_CTRL1(),
		.LPBK_IND_CTRL2(),
		.LPBK_RG_CTRL(),
		.OOBDIVCTL(),
		.OOB_PWRUP(),
		.PCI3_AUTO_REALIGN(),
		.PCI3_PIPE_RX_ELECIDLE(),
		.PCI3_RX_ASYNC_EBUF_BYPASS(),
		.PCI3_RX_ELECIDLE_EI2_ENABLE(),
		.PCI3_RX_ELECIDLE_H2L_COUNT(),
		.PCI3_RX_ELECIDLE_H2L_DISABLE(),
		.PCI3_RX_ELECIDLE_HI_COUNT(),
		.PCI3_RX_ELECIDLE_LP4_DISABLE(),
		.PCI3_RX_FIFO_DISABLE(),
		.PCIE3_CLK_COR_EMPTY_THRSH(),
		.PCIE3_CLK_COR_FULL_THRSH(),
		.PCIE3_CLK_COR_MAX_LAT(),
		.PCIE3_CLK_COR_MIN_LAT(),
		.PCIE3_CLK_COR_THRSH_TIMER(),
		.PCIE_64B_DYN_CLKSW_DIS(),
		.PCIE_BUFG_DIV_CTRL(),
		.PCIE_GEN4_64BIT_INT_EN(),
		.PCIE_PLL_SEL_MODE_GEN12(),
		.PCIE_PLL_SEL_MODE_GEN3(),
		.PCIE_PLL_SEL_MODE_GEN4(),
		.PCIE_RXPCS_CFG_GEN3(),
		.PCIE_RXPMA_CFG(),
		.PCIE_TXPCS_CFG_GEN3(),
		.PCIE_TXPMA_CFG(),
		.PCS_PCIE_EN(),
		.PCS_RSVD0(),
		.PD_TRANS_TIME_FROM_P2(),
		.PD_TRANS_TIME_NONE_P2(),
		.PD_TRANS_TIME_TO_P2(),
		.PREIQ_FREQ_BST(),
		.RATE_SW_USE_DRP(),
		.RCLK_SIPO_DLY_ENB(),
		.RCLK_SIPO_INV_EN(),
		.RTX_BUF_CML_CTRL(),
		.RTX_BUF_TERM_CTRL(),
		.RXBUFRESET_TIME(),
		.RXBUF_ADDR_MODE(),
		.RXBUF_EIDLE_HI_CNT(),
		.RXBUF_EIDLE_LO_CNT(),
		.RXBUF_EN(),
		.RXBUF_RESET_ON_CB_CHANGE(),
		.RXBUF_RESET_ON_COMMAALIGN(),
		.RXBUF_RESET_ON_EIDLE(),
		.RXBUF_RESET_ON_RATE_CHANGE(),
		.RXBUF_THRESH_OVFLW(),
		.RXBUF_THRESH_OVRD(),
		.RXBUF_THRESH_UNDFLW(),
		.RXCDRFREQRESET_TIME(),
		.RXCDRPHRESET_TIME(),
		.RXCDR_CFG0(),
		.RXCDR_CFG0_GEN3(),
		.RXCDR_CFG1(),
		.RXCDR_CFG1_GEN3(),
		.RXCDR_CFG2(),
		.RXCDR_CFG2_GEN2(),
		.RXCDR_CFG2_GEN3(),
		.RXCDR_CFG2_GEN4(),
		.RXCDR_CFG3(),
		.RXCDR_CFG3_GEN2(),
		.RXCDR_CFG3_GEN3(),
		.RXCDR_CFG3_GEN4(),
		.RXCDR_CFG4(),
		.RXCDR_CFG4_GEN3(),
		.RXCDR_CFG5(),
		.RXCDR_CFG5_GEN3(),
		.RXCDR_FR_RESET_ON_EIDLE(),
		.RXCDR_HOLD_DURING_EIDLE(),
		.RXCDR_LOCK_CFG0(),
		.RXCDR_LOCK_CFG1(),
		.RXCDR_LOCK_CFG2(),
		.RXCDR_LOCK_CFG3(),
		.RXCDR_LOCK_CFG4(),
		.RXCDR_PH_RESET_ON_EIDLE(),
		.RXCFOK_CFG0(),
		.RXCFOK_CFG1(),
		.RXCFOK_CFG2(),
		.RXCKCAL1_IQ_LOOP_RST_CFG(),
		.RXCKCAL1_I_LOOP_RST_CFG(),
		.RXCKCAL1_Q_LOOP_RST_CFG(),
		.RXCKCAL2_DX_LOOP_RST_CFG(),
		.RXCKCAL2_D_LOOP_RST_CFG(),
		.RXCKCAL2_S_LOOP_RST_CFG(),
		.RXCKCAL2_X_LOOP_RST_CFG(),
		.RXDFELPMRESET_TIME(),
		.RXDFELPM_KL_CFG0(),
		.RXDFELPM_KL_CFG1(),
		.RXDFELPM_KL_CFG2(),
		.RXDFE_CFG0(),
		.RXDFE_CFG1(),
		.RXDFE_GC_CFG0(),
		.RXDFE_GC_CFG1(),
		.RXDFE_GC_CFG2(),
		.RXDFE_H2_CFG0(),
		.RXDFE_H2_CFG1(),
		.RXDFE_H3_CFG0(),
		.RXDFE_H3_CFG1(),
		.RXDFE_H4_CFG0(),
		.RXDFE_H4_CFG1(),
		.RXDFE_H5_CFG0(),
		.RXDFE_H5_CFG1(),
		.RXDFE_H6_CFG0(),
		.RXDFE_H6_CFG1(),
		.RXDFE_H7_CFG0(),
		.RXDFE_H7_CFG1(),
		.RXDFE_H8_CFG0(),
		.RXDFE_H8_CFG1(),
		.RXDFE_H9_CFG0(),
		.RXDFE_H9_CFG1(),
		.RXDFE_HA_CFG0(),
		.RXDFE_HA_CFG1(),
		.RXDFE_HB_CFG0(),
		.RXDFE_HB_CFG1(),
		.RXDFE_HC_CFG0(),
		.RXDFE_HC_CFG1(),
		.RXDFE_HD_CFG0(),
		.RXDFE_HD_CFG1(),
		.RXDFE_HE_CFG0(),
		.RXDFE_HE_CFG1(),
		.RXDFE_HF_CFG0(),
		.RXDFE_HF_CFG1(),
		.RXDFE_KH_CFG0(),
		.RXDFE_KH_CFG1(),
		.RXDFE_KH_CFG2(),
		.RXDFE_KH_CFG3(),
		.RXDFE_OS_CFG0(),
		.RXDFE_OS_CFG1(),
		.RXDFE_UT_CFG0(),
		.RXDFE_UT_CFG1(),
		.RXDFE_UT_CFG2(),
		.RXDFE_VP_CFG0(),
		.RXDFE_VP_CFG1(),
		.RXDLY_CFG(),
		.RXDLY_LCFG(),
		.RXELECIDLE_CFG(),
		.RXGBOX_FIFO_INIT_RD_ADDR(),
		.RXGEARBOX_EN(),
		.RXISCANRESET_TIME(),
		.RXLPM_CFG(),
		.RXLPM_GC_CFG(),
		.RXLPM_KH_CFG0(),
		.RXLPM_KH_CFG1(),
		.RXLPM_OS_CFG0(),
		.RXLPM_OS_CFG1(),
		.RXOOB_CFG(),
		.RXOOB_CLK_CFG(),
		.RXOSCALRESET_TIME(),
		.RXOUT_DIV(),
		.RXPCSRESET_TIME(),
		.RXPHBEACON_CFG(),
		.RXPHDLY_CFG(),
		.RXPHSAMP_CFG(),
		.RXPHSLIP_CFG(),
		.RXPH_MONITOR_SEL(),
		.RXPI_CFG0(),
		.RXPI_CFG1(),
		.RXPMACLK_SEL(),
		.RXPMARESET_TIME(),
		.RXPRBS_ERR_LOOPBACK(),
		.RXPRBS_LINKACQ_CNT(),
		.RXREFCLKDIV2_SEL(),
		.RXSLIDE_AUTO_WAIT(),
		.RXSLIDE_MODE(),
		.RXSYNC_MULTILANE(),
		.RXSYNC_OVRD(),
		.RXSYNC_SKIP_DA(),
		.RX_AFE_CM_EN(),
		.RX_BIAS_CFG0(),
		.RX_BUFFER_CFG(),
		.RX_CAPFF_SARC_ENB(),
		.RX_CLK25_DIV(),
		.RX_CLKMUX_EN(),
		.RX_CLK_SLIP_OVRD(),
		.RX_CM_BUF_CFG(),
		.RX_CM_BUF_PD(),
		.RX_CM_SEL(),
		.RX_CM_TRIM(),
		.RX_CTLE_PWR_SAVING(),
		.RX_CTLE_RES_CTRL(),
		.RX_DATA_WIDTH(),
		.RX_DDI_SEL(),
		.RX_DEFER_RESET_BUF_EN(),
		.RX_DEGEN_CTRL(),
		.RX_DFELPM_CFG0(),
		.RX_DFELPM_CFG1(),
		.RX_DFELPM_KLKH_AGC_STUP_EN(),
		.RX_DFE_AGC_CFG1(),
		.RX_DFE_KL_LPM_KH_CFG0(),
		.RX_DFE_KL_LPM_KH_CFG1(),
		.RX_DFE_KL_LPM_KL_CFG0(),
		.RX_DFE_KL_LPM_KL_CFG1(),
		.RX_DFE_LPM_HOLD_DURING_EIDLE(),
		.RX_DISPERR_SEQ_MATCH(),
		.RX_DIVRESET_TIME(),
		.RX_EN_CTLE_RCAL_B(),
		.RX_EN_SUM_RCAL_B(),
		.RX_EYESCAN_VS_CODE(),
		.RX_EYESCAN_VS_NEG_DIR(),
		.RX_EYESCAN_VS_RANGE(),
		.RX_EYESCAN_VS_UT_SIGN(),
		.RX_FABINT_USRCLK_FLOP(),
		.RX_I2V_FILTER_EN(),
		.RX_INT_DATAWIDTH(),
		.RX_PMA_POWER_SAVE(),
		.RX_PMA_RSV0(),
		.RX_PROGDIV_CFG(),
		.RX_PROGDIV_RATE(),
		.RX_RESLOAD_CTRL(),
		.RX_RESLOAD_OVRD(),
		.RX_SAMPLE_PERIOD(),
		.RX_SIG_VALID_DLY(),
		.RX_SUM_DEGEN_AVTT_OVERITE(),
		.RX_SUM_DFETAPREP_EN(),
		.RX_SUM_IREF_TUNE(),
		.RX_SUM_PWR_SAVING(),
		.RX_SUM_RES_CTRL(),
		.RX_SUM_VCMTUNE(),
		.RX_SUM_VCM_BIAS_TUNE_EN(),
		.RX_SUM_VCM_OVWR(),
		.RX_SUM_VREF_TUNE(),
		.RX_TUNE_AFE_OS(),
		.RX_VREG_CTRL(),
		.RX_VREG_PDB(),
		.RX_WIDEMODE_CDR(),
		.RX_WIDEMODE_CDR_GEN3(),
		.RX_WIDEMODE_CDR_GEN4(),
		.RX_XCLK_SEL(),
		.RX_XMODE_SEL(),
		.SAMPLE_CLK_PHASE(),
		.SAS_12G_MODE(),
		.SATA_BURST_SEQ_LEN(),
		.SATA_BURST_VAL(),
		.SATA_CPLL_CFG(),
		.SATA_EIDLE_VAL(),
		.SHOW_REALIGN_COMMA(),
		.SIM_MODE(),
		.SIM_RECEIVER_DETECT_PASS(),
		.SIM_RESET_SPEEDUP(),
		.SIM_TX_EIDLE_DRIVE_LEVEL(),
		.SIM_DEVICE(),
		.SRSTMODE(),
		.TAPDLY_SET_TX(),
		.TERM_RCAL_CFG(),
		.TERM_RCAL_OVRD(),
		.TRANS_TIME_RATE(),
		.TST_RSV0(),
		.TST_RSV1(),
		.TXBUF_EN(),
		.TXBUF_RESET_ON_RATE_CHANGE(),
		.TXDLY_CFG(),
		.TXDLY_LCFG(),
		.TXDRV_FREQBAND(),
		.TXFE_CFG0(),
		.TXFE_CFG1(),
		.TXFE_CFG2(),
		.TXFE_CFG3(),
		.TXFIFO_ADDR_CFG(),
		.TXGBOX_FIFO_INIT_RD_ADDR(),
		.TXGEARBOX_EN(),
		.TXOUT_DIV(),
		.TXPCSRESET_TIME(),
		.TXPHDLY_CFG0(),
		.TXPHDLY_CFG1(),
		.TXPH_CFG(),
		.TXPH_CFG2(),
		.TXPH_MONITOR_SEL(),
		.TXPI_CFG0(),
		.TXPI_CFG1(),
		.TXPI_GRAY_SEL(),
		.TXPI_INVSTROBE_SEL(),
		.TXPI_PPM(),
		.TXPI_PPM_CFG(),
		.TXPI_SYNFREQ_PPM(),
		.TXPMARESET_TIME(),
		.TXREFCLKDIV2_SEL(),
		.TXSWBST_BST(),
		.TXSWBST_EN(),
		.TXSWBST_MAG(),
		.TXSYNC_MULTILANE(),
		.TXSYNC_OVRD(),
		.TXSYNC_SKIP_DA(),
		.TX_CLK25_DIV(),
		.TX_CLKMUX_EN(),
		.TX_DATA_WIDTH(),
		.TX_DCC_LOOP_RST_CFG(),
		.TX_DEEMPH0(),
		.TX_DEEMPH1(),
		.TX_DEEMPH2(),
		.TX_DEEMPH3(),
		.TX_DIVRESET_TIME(),
		.TX_DRIVE_MODE(),
		.TX_EIDLE_ASSERT_DELAY(),
		.TX_EIDLE_DEASSERT_DELAY(),
		.TX_FABINT_USRCLK_FLOP(),
		.TX_FIFO_BYP_EN(),
		.TX_IDLE_DATA_ZERO(),
		.TX_INT_DATAWIDTH(),
		.TX_LOOPBACK_DRIVE_HIZ(),
		.TX_MAINCURSOR_SEL(),
		.TX_MARGIN_FULL_0(),
		.TX_MARGIN_FULL_1(),
		.TX_MARGIN_FULL_2(),
		.TX_MARGIN_FULL_3(),
		.TX_MARGIN_FULL_4(),
		.TX_MARGIN_LOW_0(),
		.TX_MARGIN_LOW_1(),
		.TX_MARGIN_LOW_2(),
		.TX_MARGIN_LOW_3(),
		.TX_MARGIN_LOW_4(),
		.TX_PHICAL_CFG0(),
		.TX_PHICAL_CFG1(),
		.TX_PI_BIASSET(),
		.TX_PMADATA_OPT(),
		.TX_PMA_POWER_SAVE(),
		.TX_PMA_RSV0(),
		.TX_PMA_RSV1(),
		.TX_PROGCLK_SEL(),
		.TX_PROGDIV_CFG(),
		.TX_PROGDIV_RATE(),
		.TX_RXDETECT_CFG(),
		.TX_RXDETECT_REF(),
		.TX_SAMPLE_PERIOD(),
		.TX_SW_MEAS(),
		.TX_VREG_CTRL(),
		.TX_VREG_PDB(),
		.TX_VREG_VREFSEL(),
		.TX_XCLK_SEL(),
		.USB_BOTH_BURST_IDLE(),
		.USB_BURSTMAX_U3WAKE(),
		.USB_BURSTMIN_U3WAKE(),
		.USB_CLK_COR_EQ_EN(),
		.USB_EXT_CNTL(),
		.USB_IDLEMAX_POLLING(),
		.USB_IDLEMIN_POLLING(),
		.USB_LFPSPING_BURST(),
		.USB_LFPSPOLLING_BURST(),
		.USB_LFPSPOLLING_IDLE_MS(),
		.USB_LFPSU1EXIT_BURST(),
		.USB_LFPSU2LPEXIT_BURST_MS(),
		.USB_LFPSU3WAKE_BURST_MS(),
		.USB_LFPS_TPERIOD(),
		.USB_LFPS_TPERIOD_ACCURATE(),
		.USB_MODE(),
		.USB_PCIE_ERR_REP_DIS(),
		.USB_PING_SATA_MAX_INIT(),
		.USB_PING_SATA_MIN_INIT(),
		.USB_POLL_SATA_MAX_BURST(),
		.USB_POLL_SATA_MIN_BURST(),
		.USB_RAW_ELEC(),
		.USB_RXIDLE_P0_CTRL(),
		.USB_TXIDLE_TUNE_ENABLE(),
		.USB_U1_SATA_MAX_WAKE(),
		.USB_U1_SATA_MIN_WAKE(),
		.USB_U2_SAS_MAX_COM(),
		.USB_U2_SAS_MIN_COM(),
		.USE_PCS_CLK_PHASE_SEL(),
		.Y_ALL_MODE()
	) channel (

		//Top level ports
		.GTYRXP(),
		.GTYRXN(),

		.GTYTXP(),
		.GTYTXN(),

		//Data
		.TXDATA(),
		.TXDATAEXTENDRSVD(),

		.RXDATA(),
		.RXDATAEXTENDRSVD(),
		.RXDATAVALID(),
		.RXHEADER(),
		.RXHEADERVALID(),

		//Idle, power down, and loopback controls
		.RXELECIDLEMODE(),
		.RXELECIDLE(),
		.RXPD(),
		.LOOPBACK(),

		//TX driver control
		.TXDEEMPH(),
		.TXDIFFCTRL(),
		.TXELECIDLE(),
		.TXINHIBIT(),
		.TXMAINCURSOR(),
		.TXMARGIN(),
		.TXPD(),
		.TXPDELECIDLEMODE(),
		.TXPOLARITY(),
		.TXPOSTCURSOR(),
		.TXPRECURSOR(),
		.TXSWING(),

		//RX PHY controls
		.RXPOLARITY(),
		.RXTERMINATION(),

		//Reference clocks
		.GTGREFCLK(),
		.GTNORTHREFCLK0(),
		.GTNORTHREFCLK1(),
		.GTREFCLK0(),
		.GTREFCLK1(),
		.GTSOUTHREFCLK0(),
		.GTSOUTHREFCLK1(),

		//Input clocks
		.RXLATCLK(),
		.RXUSERRDY(),
		.RXUSRCLK(),
		.RXUSRCLK2(),
		.SIGVALIDCLK(),
		.TXLATCLK(),
		.TXPHDLYTSTCLK(),
		.TXUSERRDY(),
		.TXUSRCLK(),
		.TXUSRCLK2(),

		//Output clocks
		.RXOUTCLKSEL(),
		.RXPLLCLKSEL(),
		.RXSLIPOUTCLK(),
		.RXSYSCLKSEL(),
		.TXOUTCLKSEL(),
		.TXPLLCLKSEL(),
		.TXSYSCLKSEL(),
		.RXOUTCLK(),
		.RXOUTCLKFABRIC(),
		.RXOUTCLKPCS(),
		.RXRECCLKOUT(),
		.TXOUTCLK(),
		.TXOUTCLKFABRIC(),
		.TXOUTCLKPCS(),

		//Clock outputs or something?
		.BUFGTCE(),
		.BUFGTCEMASK(),
		.BUFGTDIV(),

		//Clocks and status inputs from QPLL
		.QPLL0CLK(),
		.QPLL0FREQLOCK(),
		.QPLL0REFCLK(),
		.QPLL1CLK(),
		.QPLL1FREQLOCK(),
		.QPLL1REFCLK(),

		//CPLL status outputs
		.CPLLFBCLKLOST(),
		.CPLLLOCK(),
		.CPLLREFCLKLOST(),

		//Sub-rate control
		.RXRATE(),
		.RXRATEMODE(),
		.TXRATE(),
		.TXRATEMODE(),
		.RXRATEDONE(),
		.TXRATEDONE(),

		//Resets
		.GTRXRESET(),
		.GTRXRESETSEL(),
		.GTTXRESET(),
		.GTTXRESETSEL(),
		.RESETOVRD(),
		.RXBUFRESET(),
		.RXCDRFREQRESET(),
		.RXCDRRESET(),
		.RXCKCALRESET(),
		.RXDFELPMRESET(),
		.RXDLYSRESET(),
		.RXOOBRESET(),
		.RXOSCALRESET(),
		.RXPCSRESET(),
		.RXPHDLYRESET(),
		.RXPMARESET(),
		.RXPROGDIVRESET(),
		.TXDCCRESET(),
		.TXDLYSRESET(),
		.TXLFPSTRESET(),
		.TXPCSRESET(),
		.TXPHDLYRESET(),
		.TXPMARESET(),
		.TXPROGDIVRESET(),
		.BUFGTRESET(),
		.BUFGTRSTMASK(),

		.RXDLYSRESETDONE(),
		.RXPMARESETDONE(),
		.RXPRGDIVRESETDONE(),
		.RXRESETDONE(),
		.TXDLYSRESETDONE(),
		.TXPMARESETDONE(),
		.TXPRGDIVRESETDONE(),
		.TXRESETDONE(),

		//PRBS generator and checker
		.RXPRBSCNTRESET(),
		.RXPRBSSEL(),
		.TXPRBSFORCEERR(),
		.TXPRBSSEL(),
		.RXPRBSERR(),
		.RXPRBSLOCKED(),

		//RX 8B10B decoder and comma aligner
		.RX8B10BEN(),
		.RXCOMMADETEN(),
		.RXMCOMMAALIGNEN(),
		.RXPCOMMAALIGNEN(),
		.RXBYTEISALIGNED(),
		.RXBYTEREALIGN(),
		.RXCOMMADET(),

		//RX CDR
		.RXCDRHOLD(),
		.RXCDROVRDEN(),
		.RXCDRLOCK(),
		.RXCDRPHDONE(),

		//RX channel bonding
		.RXCHBONDEN(),
		.RXCHBONDI(),
		.RXCHBONDLEVEL(),
		.RXCHBONDMASTER(),
		.RXCHBONDSLAVE(),
		.RXCHANBONDSEQ(),
		.RXCHANISALIGNED(),
		.RXCHANREALIGN(),
		.RXCHBONDO(),

		//RX CTLE
		.RXLPMEN(),
		.RXLPMGCHOLD(),
		.RXLPMGCOVRDEN(),
		.RXLPMHFHOLD(),
		.RXLPMHFOVRDEN(),
		.RXLPMLFHOLD(),
		.RXLPMLFKLOVRDEN(),
		.RXLPMOSHOLD(),
		.RXLPMOSOVRDEN(),

		//RX DFE
		.RXDFEAGCHOLD(),
		.RXDFEAGCOVRDEN(),
		.RXDFECFOKFCNUM(),
		.RXDFECFOKFEN(),
		.RXDFECFOKFPULSE(),
		.RXDFECFOKHOLD(),
		.RXDFECFOKOVREN(),
		.RXDFEKHHOLD(),
		.RXDFEKHOVRDEN(),
		.RXDFELFHOLD(),
		.RXDFELFOVRDEN(),
		.RXDFETAP2HOLD(),
		.RXDFETAP2OVRDEN(),
		.RXDFETAP3HOLD(),
		.RXDFETAP3OVRDEN(),
		.RXDFETAP4HOLD(),
		.RXDFETAP4OVRDEN(),
		.RXDFETAP5HOLD(),
		.RXDFETAP5OVRDEN(),
		.RXDFETAP6HOLD(),
		.RXDFETAP6OVRDEN(),
		.RXDFETAP7HOLD(),
		.RXDFETAP7OVRDEN(),
		.RXDFETAP8HOLD(),
		.RXDFETAP8OVRDEN(),
		.RXDFETAP9HOLD(),
		.RXDFETAP9OVRDEN(),
		.RXDFETAP10HOLD(),
		.RXDFETAP10OVRDEN(),
		.RXDFETAP11HOLD(),
		.RXDFETAP11OVRDEN(),
		.RXDFETAP12HOLD(),
		.RXDFETAP12OVRDEN(),
		.RXDFETAP13HOLD(),
		.RXDFETAP13OVRDEN(),
		.RXDFETAP14HOLD(),
		.RXDFETAP14OVRDEN(),
		.RXDFETAP15HOLD(),
		.RXDFETAP15OVRDEN(),
		.RXDFEUTHOLD(),
		.RXDFEUTOVRDEN(),
		.RXDFEVPHOLD(),
		.RXDFEVPOVRDEN(),
		.RXDFEXYDEN(),

		//RX delay
		.RXDLYBYPASS(),
		.RXDLYEN(),
		.RXDLYOVRDEN(),

		//RX phase aligner
		.RXPHALIGN(),
		.RXPHALIGNEN(),
		.RXPHDLYPD(),
		.RXPHALIGNDONE(),
		.RXPHALIGNERR(),

		//TX 8B/10B coder
		.TX8B10BBYPASS(),
		.TX8B10BEN(),

		//TX gearbox
		.TXHEADER(),
		.TXSEQUENCE(),

		//SATA/SAS (not used)
		.TXCOMINIT(),
		.TXCOMSAS(),
		.TXCOMWAKE(),
		.TXCOMFINISH(),
		.RXCOMINITDET(),
		.RXCOMSASDET(),
		.RXCOMWAKEDET(),

		//TX delay
		.TXDLYBYPASS(),
		.TXDLYEN(),
		.TXDLYHOLD(),
		.TXDLYOVRDEN(),
		.TXDLYUPDOWN(),

		//TX phase aligner
		.TXPHALIGN(),
		.TXPHALIGNEN(),
		.TXPHDLYPD(),
		.TXPHINIT(),
		.TXPHOVRDEN(),

		//TX interpolator
		.TXPIPPMEN(),
		.TXPIPPMOVRDEN(),
		.TXPIPPMPD(),
		.TXPIPPMSEL(),
		.TXPIPPMSTEPSIZE(),

		//TODO
		.TXSYNCDONE(),
		.TXSYNCOUT(),
		.RXSLIDERDY(),
		.RXSLIPDONE(),
		.RXSLIPOUTCLKRDY(),
		.RXSLIPPMARDY(),
		.RXSTARTOFSEQ(),
		.RXSTATUS(),
		.RXSYNCDONE(),
		.RXSYNCOUT(),
		.RXVALID(),
		.TXBUFSTATUS(),
		.RXLFPSTRESETDET(),
		.RXLFPSU2LPEXITDET(),
		.RXLFPSU3WAKEDET(),
		.RXMONITOROUT(),
		.RXOSINTDONE(),
		.RXOSINTSTARTED(),
		.RXOSINTSTROBEDONE(),
		.RXOSINTSTROBESTARTED(),
		.RXCTRL0(),
		.RXCTRL1(),
		.RXCTRL2(),
		.RXCTRL3(),
		.RXCKCALDONE(),
		.RXCLKCORCNT(),
		.RXBUFSTATUS(),
		.PHYSTATUS(),
		.PINRSRVDAS(),
		.POWERPRESENT(),
		.RESETEXCEPTION(),
		.GTPOWERGOOD(),
		.GTREFCLKMONITOR(),
		.EYESCANDATAERROR(),
		.DMONITOROUT(),
		.DMONITOROUTCLK(),
		.TXSYNCALLIN(),
		.TXSYNCIN(),
		.TXSYNCMODE(),
		.TXPISOPD(),
		.TXMUXDCDEXHOLD(),
		.TXMUXDCDORWREN(),
		.TXONESZEROS(),
		.TXLFPSU2LPEXIT(),
		.TXLFPSU3WAKE(),
		.TXDETECTRX(),
		.TXDCCFORCESTART(),
		.TXCTRL0(),
		.TXCTRL1(),
		.TXCTRL2(),
		.TSTIN(),
		.RXSYNCALLIN(),
		.RXSYNCIN(),
		.RXSYNCMODE(),
		.RXSLIDE(),
		.RXSLIPPMA(),
		.RXMONITORSEL(),
		.RXEQTRAINING(),
		.RXGEARBOXSLIP(),
		.RXCKCALSTART(),
		.RXAFECFOKEN(),
		.CDRSTEPDIR(),
		.CDRSTEPSQ(),
		.CDRSTEPSX(),
		.CFGRESET(),
		.CLKRSVD0(),
		.CLKRSVD1(),
		.CPLLFREQLOCK(),
		.CPLLLOCKDETCLK(),
		.CPLLLOCKEN(),
		.CPLLPD(),
		.CPLLREFCLKSEL(),
		.CPLLRESET(),
		.DMONFIFORESET(),
		.DMONITORCLK(),
		.EYESCANRESET(),
		.EYESCANTRIGGER(),
		.FREQOS(),
		.GTRSVD(),
		.INCPCTRL(),
		.RXOSHOLD(),
		.RXOSOVRDEN(),
		.TXDCCDONE(),
		.TXPHALIGNDONE(),
		.TXPHINITDONE(),

		//PCIe mode, ignore for now
		.PCIEEQRXEQADAPTDONE(),
		.PCIERSTIDLE(),
		.PCIERSTTXSYNCSTART(),
		.PCIEUSERRATEDONE(),
		.PCSRSVDIN(),
		.PCIERATEGEN3(),
		.PCIERATEIDLE(),
		.PCIERATEQPLLPD(),
		.PCIERATEQPLLRESET(),
		.PCIESYNCTXSYNCDONE(),
		.PCIEUSERGEN3RDY(),
		.PCIEUSERPHYSTATUSRST(),
		.PCIEUSERRATESTART(),
		.PCSRSVDOUT(),

		//DRP (bridged to APB)
		.DRPADDR(),
		.DRPCLK(),
		.DRPDI(),
		.DRPEN(),
		.DRPRST(),
		.DRPWE(),
		.DRPDO(),
		.DRPRDY()

		//Reserved ports, ignore or tie off.
	);

endmodule
